<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" id="terminal" baseProfile="full" viewBox="0 0 500 430" width="550" version="1.1">
    <defs>
        <termtosvg:template_settings xmlns:termtosvg="https://github.com/nbedos/termtosvg">
            <termtosvg:screen_geometry columns="95" rows="21" />
            <termtosvg:animation type="css" />
        </termtosvg:template_settings>
        <style type="text/css" id="generated-style">
            <![CDATA[#screen {
                font-family: 'DejaVu Sans Mono', monospace;
                font-style: normal;
                font-size: 14px;
            }

        text {
            dominant-baseline: text-before-edge;
            white-space: pre;
        }
    
            :root {
                --animation-duration: 14558ms;
            }

            @keyframes roll {
                0.000%{transform:translateY(0px)}
3.400%{transform:translateY(-374px)}
4.767%{transform:translateY(-748px)}
7.302%{transform:translateY(-1122px)}
9.933%{transform:translateY(-1496px)}
12.357%{transform:translateY(-1870px)}
14.226%{transform:translateY(-2244px)}
17.578%{transform:translateY(-2618px)}
21.239%{transform:translateY(-2992px)}
21.658%{transform:translateY(-3366px)}
24.605%{transform:translateY(-3740px)}
27.627%{transform:translateY(-4114px)}
29.771%{transform:translateY(-4488px)}
31.529%{transform:translateY(-4862px)}
34.277%{transform:translateY(-5236px)}
36.585%{transform:translateY(-5610px)}
39.607%{transform:translateY(-5984px)}
41.256%{transform:translateY(-6358px)}
43.179%{transform:translateY(-6732px)}
44.333%{transform:translateY(-7106px)}
47.685%{transform:translateY(-7480px)}
51.436%{transform:translateY(-7854px)}
51.889%{transform:translateY(-8228px)}
59.658%{transform:translateY(-8602px)}
62.241%{transform:translateY(-8976px)}
64.885%{transform:translateY(-9350px)}
67.406%{transform:translateY(-9724px)}
68.347%{transform:translateY(-10098px)}
70.985%{transform:translateY(-10472px)}
77.469%{transform:translateY(-10846px)}
81.124%{transform:translateY(-11220px)}
81.536%{transform:translateY(-11594px)}
85.046%{transform:translateY(-11968px)}
86.090%{transform:translateY(-12342px)}
89.442%{transform:translateY(-12716px)}
90.267%{transform:translateY(-13090px)}
93.014%{transform:translateY(-13464px)}
93.131%{transform:translateY(-13838px)}
100.000%{transform:translateY(-13838px)}
            }

            #screen_view {
                animation-duration: 14558ms;
                animation-iteration-count:infinite;
                animation-name:roll;
                animation-timing-function: steps(1,end);
                animation-fill-mode: forwards;
            }
        ]]>
        </style>
        <style type="text/css" id="user-style">
            /* The colors defined below are the default 16 colors used for rendering text of the terminal. Adjust
               them as needed.
               gjm8 color theme (source: https://terminal.sexy/) */
            .foreground {fill: #00FF00}
            .background {fill: #000000}
            .color0 {fill: #272822}
            .color1 {fill: #f92672}
            .green {fill: #00FF00}
            .color3 {fill: #f4bf75}
            .color4 {fill: #66d9ef}
            .purple {fill: #00FF00}
            .color6 {fill: #00FF00}
            .color7 {fill: #f8f8f2}
            .color8 {fill: #75715e}
            .color9 {fill: #fd971f}
            .color10 {fill: #00FF00}
            .color11 {fill: #49483e}
            .color12 {fill: #00FF00}
            .color13 {fill: #f5f4f1}
            .orange {fill: #00FF00}
            .color15 {fill: #f9f8f5}
        </style>
    </defs>
    <rect id="terminalui" class="background" width="100%" height="100%" ry="4.5826941" />
    <circle cx="24" cy="23" r="7" fill="#f92672" />
    <circle cx="44" cy="23" r="7" fill="#f4bf75" />
    <circle cx="64" cy="23" r="7" fill="#a6e22e" />
    <svg id="screen" width="760" height="357" x="23" y="50" viewBox="0 0 760 357" preserveAspectRatio="xMidYMin slice">
        <rect class="background" height="100%" width="100%" x="0" y="0" />
        <defs>
            <g id="g1">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="16" class="foreground">$ </text>
                <text x="160" textLength="8" class="background"></text>
            </g>
            <g id="g2">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="24" class="foreground">$ w</text>
                <text x="168" textLength="8" class="background"></text>
            </g>
            <g id="g3">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="32" class="foreground">$ wh</text>
                <text x="176" textLength="8" class="background"></text>
            </g>
            <g id="g4">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="40" class="foreground">$ who</text>
                <text x="184" textLength="8" class="background"></text>
            </g>
            <g id="g5">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="48" class="foreground">$ whoa</text>
                <text x="192" textLength="8" class="background"></text>
            </g>
            <g id="g6">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="56" class="foreground">$ whoam</text>
                <text x="200" textLength="8" class="background"></text>
            </g>
            <g id="g7">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="64" class="foreground">$ whoami</text>
                <text x="208" textLength="8" class="background"></text>
            </g>
            <g id="g8">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="64" class="foreground">$ whoami</text>
            </g>
            <g id="g9">
                <text x="0" textLength="8" class="background"></text>
            </g>
            <g id="g10">
                <text x="0" textLength="104" class="color6">Less</text>
            </g>
            <g id="g11">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="24" class="foreground">$ g</text>
                <text x="168" textLength="8" class="background"></text>
            </g>
            <g id="g12">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="32" class="foreground">$ gi</text>
                <text x="176" textLength="8" class="background"></text>
            </g>
            <g id="g13">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="40" class="foreground">$ git</text>
                <text x="184" textLength="8" class="background"></text>
            </g>
            <g id="g14">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="48" class="foreground">$ git </text>
                <text x="192" textLength="8" class="background"></text>
            </g>
            <g id="g15">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="56" class="foreground">$ git s</text>
                <text x="200" textLength="8" class="background"></text>
            </g>
            <g id="g16">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="64" class="foreground">$ git st</text>
                <text x="208" textLength="8" class="background"></text>
            </g>
            <g id="g17">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="72" class="foreground">$ git sta</text>
                <text x="216" textLength="8" class="background"></text>
            </g>
            <g id="g18">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="80" class="foreground">$ git stat</text>
                <text x="224" textLength="8" class="background"></text>
            </g>
            <g id="g19">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="88" class="foreground">$ git statu</text>
                <text x="232" textLength="8" class="background"></text>
            </g>
            <g id="g20">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="96" class="foreground">$ git status</text>
                <text x="240" textLength="8" class="background"></text>
            </g>
            <g id="g21">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="96" class="foreground">$ git status</text>
            </g>
            <g id="g22">
                <text x="0" textLength="240" font-style="italic" class="foreground">        GitHub Status         </text>
            </g>
            <g id="g23">
                <text x="0" textLength="240" class="foreground">&#9556;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9572;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9559;</text>
            </g>
            <g id="g24">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" font-weight="bold" class="orange"> Title         </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" font-weight="bold" class="orange"> Count      </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g25">
                <text x="0" textLength="240" class="foreground">&#9567;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9532;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9472;&#9570;</text>
            </g>
            <g id="g26">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Stars         </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 3          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g27">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Forks         </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 2          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g28">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Commits       </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 1437        </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g29">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Followers     </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 0          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g30">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Pull Requests </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 394         </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g31">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Issues        </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 3          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g32">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Repository    </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 6          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g33">
                <text x="0" textLength="8" class="foreground">&#9553;</text>
                <text x="8" textLength="120" class="purple"> Gists         </text>
                <text x="128" textLength="8" class="foreground">&#9474;</text>
                <text x="136" textLength="96" class="green"> 0          </text>
                <text x="232" textLength="8" class="foreground">&#9553;</text>
            </g>
            <g id="g34">
                <text x="0" textLength="240" class="foreground">&#9562;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9575;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9552;&#9565;</text>
            </g>
            <g id="g35">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="24" class="foreground">$ u</text>
                <text x="168" textLength="8" class="background"></text>
            </g>
            <g id="g36">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="32" class="foreground">$ up</text>
                <text x="176" textLength="8" class="background"></text>
            </g>
            <g id="g37">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="40" class="foreground">$ upt</text>
                <text x="184" textLength="8" class="background"></text>
            </g>
            <g id="g38">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="48" class="foreground">$ upti</text>
                <text x="192" textLength="8" class="background"></text>
            </g>
            <g id="g39">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="56" class="foreground">$ uptim</text>
                <text x="200" textLength="8" class="background"></text>
            </g>
            <g id="g40">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="64" class="foreground">$ uptime</text>
                <text x="208" textLength="8" class="background"></text>
            </g>
            <g id="g41">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="64" class="foreground">$ uptime</text>
            </g>
            <g id="g42">
                <text x="0" textLength="32" font-weight="bold" class="orange">79</text>
            </g>
            <g id="g43">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="24" class="foreground">$ e</text>
                <text x="168" textLength="8" class="background"></text>
            </g>
            <g id="g44">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="32" class="foreground">$ ex</text>
                <text x="176" textLength="8" class="background"></text>
            </g>
            <g id="g45">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="40" class="foreground">$ exi</text>
                <text x="184" textLength="8" class="background"></text>
            </g>
            <g id="g46">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="48" class="foreground">$ exit</text>
                <text x="192" textLength="8" class="background"></text>
            </g>
            <g id="g47">
                <text x="0" textLength="128" font-weight="bold" class="color10">less-dev@git</text>
                <text x="128" textLength="8" class="foreground">:</text>
                <text x="136" textLength="8" font-weight="bold" class="color12">~</text>
                <text x="144" textLength="48" class="foreground">$ exit</text>
            </g>
            <g id="g48">
                <text x="0" textLength="32" class="foreground">exit</text>
            </g>
        </defs>
        <g id="screen_view">
            <g>
                <rect x="160" y="0" width="8" height="17" class="foreground" />
                <use xlink:href="#g1" y="0" />
            </g>
            <g>
                <rect x="168" y="374" width="8" height="17" class="foreground" />
                <use xlink:href="#g2" y="374" />
            </g>
            <g>
                <rect x="176" y="748" width="8" height="17" class="foreground" />
                <use xlink:href="#g3" y="748" />
            </g>
            <g>
                <rect x="184" y="1122" width="8" height="17" class="foreground" />
                <use xlink:href="#g4" y="1122" />
            </g>
            <g>
                <rect x="192" y="1496" width="8" height="17" class="foreground" />
                <use xlink:href="#g5" y="1496" />
            </g>
            <g>
                <rect x="200" y="1870" width="8" height="17" class="foreground" />
                <use xlink:href="#g6" y="1870" />
            </g>
            <g>
                <rect x="208" y="2244" width="8" height="17" class="foreground" />
                <use xlink:href="#g7" y="2244" />
            </g>
            <g>
                <use xlink:href="#g8" y="2618" />
                <rect x="0" y="2635" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="2635" />
            </g>
            <g>
                <use xlink:href="#g8" y="2992" />
                <use xlink:href="#g10" y="3009" />
                <rect x="0" y="3026" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="3026" />
            </g>
            <g>
                <use xlink:href="#g8" y="3366" />
                <use xlink:href="#g10" y="3383" />
                <rect x="160" y="3400" width="8" height="17" class="foreground" />
                <use xlink:href="#g1" y="3400" />
            </g>
            <g>
                <use xlink:href="#g8" y="3740" />
                <use xlink:href="#g10" y="3757" />
                <rect x="168" y="3774" width="8" height="17" class="foreground" />
                <use xlink:href="#g11" y="3774" />
            </g>
            <g>
                <use xlink:href="#g8" y="4114" />
                <use xlink:href="#g10" y="4131" />
                <rect x="176" y="4148" width="8" height="17" class="foreground" />
                <use xlink:href="#g12" y="4148" />
            </g>
            <g>
                <use xlink:href="#g8" y="4488" />
                <use xlink:href="#g10" y="4505" />
                <rect x="184" y="4522" width="8" height="17" class="foreground" />
                <use xlink:href="#g13" y="4522" />
            </g>
            <g>
                <use xlink:href="#g8" y="4862" />
                <use xlink:href="#g10" y="4879" />
                <rect x="192" y="4896" width="8" height="17" class="foreground" />
                <use xlink:href="#g14" y="4896" />
            </g>
            <g>
                <use xlink:href="#g8" y="5236" />
                <use xlink:href="#g10" y="5253" />
                <rect x="200" y="5270" width="8" height="17" class="foreground" />
                <use xlink:href="#g15" y="5270" />
            </g>
            <g>
                <use xlink:href="#g8" y="5610" />
                <use xlink:href="#g10" y="5627" />
                <rect x="208" y="5644" width="8" height="17" class="foreground" />
                <use xlink:href="#g16" y="5644" />
            </g>
            <g>
                <use xlink:href="#g8" y="5984" />
                <use xlink:href="#g10" y="6001" />
                <rect x="216" y="6018" width="8" height="17" class="foreground" />
                <use xlink:href="#g17" y="6018" />
            </g>
            <g>
                <use xlink:href="#g8" y="6358" />
                <use xlink:href="#g10" y="6375" />
                <rect x="224" y="6392" width="8" height="17" class="foreground" />
                <use xlink:href="#g18" y="6392" />
            </g>
            <g>
                <use xlink:href="#g8" y="6732" />
                <use xlink:href="#g10" y="6749" />
                <rect x="232" y="6766" width="8" height="17" class="foreground" />
                <use xlink:href="#g19" y="6766" />
            </g>
            <g>
                <use xlink:href="#g8" y="7106" />
                <use xlink:href="#g10" y="7123" />
                <rect x="240" y="7140" width="8" height="17" class="foreground" />
                <use xlink:href="#g20" y="7140" />
            </g>
            <g>
                <use xlink:href="#g8" y="7480" />
                <use xlink:href="#g10" y="7497" />
                <use xlink:href="#g21" y="7514" />
                <rect x="0" y="7531" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="7531" />
            </g>
            <g>
                <use xlink:href="#g8" y="7854" />
                <use xlink:href="#g10" y="7871" />
                <use xlink:href="#g21" y="7888" />
                <use xlink:href="#g22" y="7905" />
                <use xlink:href="#g23" y="7922" />
                <use xlink:href="#g24" y="7939" />
                <use xlink:href="#g25" y="7956" />
                <use xlink:href="#g26" y="7973" />
                <use xlink:href="#g27" y="7990" />
                <use xlink:href="#g28" y="8007" />
                <use xlink:href="#g29" y="8024" />
                <use xlink:href="#g30" y="8041" />
                <use xlink:href="#g31" y="8058" />
                <use xlink:href="#g32" y="8075" />
                <use xlink:href="#g33" y="8092" />
                <use xlink:href="#g34" y="8109" />
                <rect x="0" y="8126" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="8126" />
            </g>
            <g>
                <use xlink:href="#g8" y="8228" />
                <use xlink:href="#g10" y="8245" />
                <use xlink:href="#g21" y="8262" />
                <use xlink:href="#g22" y="8279" />
                <use xlink:href="#g23" y="8296" />
                <use xlink:href="#g24" y="8313" />
                <use xlink:href="#g25" y="8330" />
                <use xlink:href="#g26" y="8347" />
                <use xlink:href="#g27" y="8364" />
                <use xlink:href="#g28" y="8381" />
                <use xlink:href="#g29" y="8398" />
                <use xlink:href="#g30" y="8415" />
                <use xlink:href="#g31" y="8432" />
                <use xlink:href="#g32" y="8449" />
                <use xlink:href="#g33" y="8466" />
                <use xlink:href="#g34" y="8483" />
                <rect x="160" y="8500" width="8" height="17" class="foreground" />
                <use xlink:href="#g1" y="8500" />
            </g>
            <g>
                <use xlink:href="#g8" y="8602" />
                <use xlink:href="#g10" y="8619" />
                <use xlink:href="#g21" y="8636" />
                <use xlink:href="#g22" y="8653" />
                <use xlink:href="#g23" y="8670" />
                <use xlink:href="#g24" y="8687" />
                <use xlink:href="#g25" y="8704" />
                <use xlink:href="#g26" y="8721" />
                <use xlink:href="#g27" y="8738" />
                <use xlink:href="#g28" y="8755" />
                <use xlink:href="#g29" y="8772" />
                <use xlink:href="#g30" y="8789" />
                <use xlink:href="#g31" y="8806" />
                <use xlink:href="#g32" y="8823" />
                <use xlink:href="#g33" y="8840" />
                <use xlink:href="#g34" y="8857" />
                <rect x="168" y="8874" width="8" height="17" class="foreground" />
                <use xlink:href="#g35" y="8874" />
            </g>
            <g>
                <use xlink:href="#g8" y="8976" />
                <use xlink:href="#g10" y="8993" />
                <use xlink:href="#g21" y="9010" />
                <use xlink:href="#g22" y="9027" />
                <use xlink:href="#g23" y="9044" />
                <use xlink:href="#g24" y="9061" />
                <use xlink:href="#g25" y="9078" />
                <use xlink:href="#g26" y="9095" />
                <use xlink:href="#g27" y="9112" />
                <use xlink:href="#g28" y="9129" />
                <use xlink:href="#g29" y="9146" />
                <use xlink:href="#g30" y="9163" />
                <use xlink:href="#g31" y="9180" />
                <use xlink:href="#g32" y="9197" />
                <use xlink:href="#g33" y="9214" />
                <use xlink:href="#g34" y="9231" />
                <rect x="176" y="9248" width="8" height="17" class="foreground" />
                <use xlink:href="#g36" y="9248" />
            </g>
            <g>
                <use xlink:href="#g8" y="9350" />
                <use xlink:href="#g10" y="9367" />
                <use xlink:href="#g21" y="9384" />
                <use xlink:href="#g22" y="9401" />
                <use xlink:href="#g23" y="9418" />
                <use xlink:href="#g24" y="9435" />
                <use xlink:href="#g25" y="9452" />
                <use xlink:href="#g26" y="9469" />
                <use xlink:href="#g27" y="9486" />
                <use xlink:href="#g28" y="9503" />
                <use xlink:href="#g29" y="9520" />
                <use xlink:href="#g30" y="9537" />
                <use xlink:href="#g31" y="9554" />
                <use xlink:href="#g32" y="9571" />
                <use xlink:href="#g33" y="9588" />
                <use xlink:href="#g34" y="9605" />
                <rect x="184" y="9622" width="8" height="17" class="foreground" />
                <use xlink:href="#g37" y="9622" />
            </g>
            <g>
                <use xlink:href="#g8" y="9724" />
                <use xlink:href="#g10" y="9741" />
                <use xlink:href="#g21" y="9758" />
                <use xlink:href="#g22" y="9775" />
                <use xlink:href="#g23" y="9792" />
                <use xlink:href="#g24" y="9809" />
                <use xlink:href="#g25" y="9826" />
                <use xlink:href="#g26" y="9843" />
                <use xlink:href="#g27" y="9860" />
                <use xlink:href="#g28" y="9877" />
                <use xlink:href="#g29" y="9894" />
                <use xlink:href="#g30" y="9911" />
                <use xlink:href="#g31" y="9928" />
                <use xlink:href="#g32" y="9945" />
                <use xlink:href="#g33" y="9962" />
                <use xlink:href="#g34" y="9979" />
                <rect x="192" y="9996" width="8" height="17" class="foreground" />
                <use xlink:href="#g38" y="9996" />
            </g>
            <g>
                <use xlink:href="#g8" y="10098" />
                <use xlink:href="#g10" y="10115" />
                <use xlink:href="#g21" y="10132" />
                <use xlink:href="#g22" y="10149" />
                <use xlink:href="#g23" y="10166" />
                <use xlink:href="#g24" y="10183" />
                <use xlink:href="#g25" y="10200" />
                <use xlink:href="#g26" y="10217" />
                <use xlink:href="#g27" y="10234" />
                <use xlink:href="#g28" y="10251" />
                <use xlink:href="#g29" y="10268" />
                <use xlink:href="#g30" y="10285" />
                <use xlink:href="#g31" y="10302" />
                <use xlink:href="#g32" y="10319" />
                <use xlink:href="#g33" y="10336" />
                <use xlink:href="#g34" y="10353" />
                <rect x="200" y="10370" width="8" height="17" class="foreground" />
                <use xlink:href="#g39" y="10370" />
            </g>
            <g>
                <use xlink:href="#g8" y="10472" />
                <use xlink:href="#g10" y="10489" />
                <use xlink:href="#g21" y="10506" />
                <use xlink:href="#g22" y="10523" />
                <use xlink:href="#g23" y="10540" />
                <use xlink:href="#g24" y="10557" />
                <use xlink:href="#g25" y="10574" />
                <use xlink:href="#g26" y="10591" />
                <use xlink:href="#g27" y="10608" />
                <use xlink:href="#g28" y="10625" />
                <use xlink:href="#g29" y="10642" />
                <use xlink:href="#g30" y="10659" />
                <use xlink:href="#g31" y="10676" />
                <use xlink:href="#g32" y="10693" />
                <use xlink:href="#g33" y="10710" />
                <use xlink:href="#g34" y="10727" />
                <rect x="208" y="10744" width="8" height="17" class="foreground" />
                <use xlink:href="#g40" y="10744" />
            </g>
            <g>
                <use xlink:href="#g8" y="10846" />
                <use xlink:href="#g10" y="10863" />
                <use xlink:href="#g21" y="10880" />
                <use xlink:href="#g22" y="10897" />
                <use xlink:href="#g23" y="10914" />
                <use xlink:href="#g24" y="10931" />
                <use xlink:href="#g25" y="10948" />
                <use xlink:href="#g26" y="10965" />
                <use xlink:href="#g27" y="10982" />
                <use xlink:href="#g28" y="10999" />
                <use xlink:href="#g29" y="11016" />
                <use xlink:href="#g30" y="11033" />
                <use xlink:href="#g31" y="11050" />
                <use xlink:href="#g32" y="11067" />
                <use xlink:href="#g33" y="11084" />
                <use xlink:href="#g34" y="11101" />
                <use xlink:href="#g41" y="11118" />
                <rect x="0" y="11135" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="11135" />
            </g>
            <g>
                <use xlink:href="#g8" y="11220" />
                <use xlink:href="#g10" y="11237" />
                <use xlink:href="#g21" y="11254" />
                <use xlink:href="#g22" y="11271" />
                <use xlink:href="#g23" y="11288" />
                <use xlink:href="#g24" y="11305" />
                <use xlink:href="#g25" y="11322" />
                <use xlink:href="#g26" y="11339" />
                <use xlink:href="#g27" y="11356" />
                <use xlink:href="#g28" y="11373" />
                <use xlink:href="#g29" y="11390" />
                <use xlink:href="#g30" y="11407" />
                <use xlink:href="#g31" y="11424" />
                <use xlink:href="#g32" y="11441" />
                <use xlink:href="#g33" y="11458" />
                <use xlink:href="#g34" y="11475" />
                <use xlink:href="#g41" y="11492" />
                <use xlink:href="#g42" y="11509" />
                <rect x="0" y="11526" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="11526" />
            </g>
            <g>
                <use xlink:href="#g8" y="11594" />
                <use xlink:href="#g10" y="11611" />
                <use xlink:href="#g21" y="11628" />
                <use xlink:href="#g22" y="11645" />
                <use xlink:href="#g23" y="11662" />
                <use xlink:href="#g24" y="11679" />
                <use xlink:href="#g25" y="11696" />
                <use xlink:href="#g26" y="11713" />
                <use xlink:href="#g27" y="11730" />
                <use xlink:href="#g28" y="11747" />
                <use xlink:href="#g29" y="11764" />
                <use xlink:href="#g30" y="11781" />
                <use xlink:href="#g31" y="11798" />
                <use xlink:href="#g32" y="11815" />
                <use xlink:href="#g33" y="11832" />
                <use xlink:href="#g34" y="11849" />
                <use xlink:href="#g41" y="11866" />
                <use xlink:href="#g42" y="11883" />
                <rect x="160" y="11900" width="8" height="17" class="foreground" />
                <use xlink:href="#g1" y="11900" />
            </g>
            <g>
                <use xlink:href="#g8" y="11968" />
                <use xlink:href="#g10" y="11985" />
                <use xlink:href="#g21" y="12002" />
                <use xlink:href="#g22" y="12019" />
                <use xlink:href="#g23" y="12036" />
                <use xlink:href="#g24" y="12053" />
                <use xlink:href="#g25" y="12070" />
                <use xlink:href="#g26" y="12087" />
                <use xlink:href="#g27" y="12104" />
                <use xlink:href="#g28" y="12121" />
                <use xlink:href="#g29" y="12138" />
                <use xlink:href="#g30" y="12155" />
                <use xlink:href="#g31" y="12172" />
                <use xlink:href="#g32" y="12189" />
                <use xlink:href="#g33" y="12206" />
                <use xlink:href="#g34" y="12223" />
                <use xlink:href="#g41" y="12240" />
                <use xlink:href="#g42" y="12257" />
                <rect x="168" y="12274" width="8" height="17" class="foreground" />
                <use xlink:href="#g43" y="12274" />
            </g>
            <g>
                <use xlink:href="#g8" y="12342" />
                <use xlink:href="#g10" y="12359" />
                <use xlink:href="#g21" y="12376" />
                <use xlink:href="#g22" y="12393" />
                <use xlink:href="#g23" y="12410" />
                <use xlink:href="#g24" y="12427" />
                <use xlink:href="#g25" y="12444" />
                <use xlink:href="#g26" y="12461" />
                <use xlink:href="#g27" y="12478" />
                <use xlink:href="#g28" y="12495" />
                <use xlink:href="#g29" y="12512" />
                <use xlink:href="#g30" y="12529" />
                <use xlink:href="#g31" y="12546" />
                <use xlink:href="#g32" y="12563" />
                <use xlink:href="#g33" y="12580" />
                <use xlink:href="#g34" y="12597" />
                <use xlink:href="#g41" y="12614" />
                <use xlink:href="#g42" y="12631" />
                <rect x="176" y="12648" width="8" height="17" class="foreground" />
                <use xlink:href="#g44" y="12648" />
            </g>
            <g>
                <use xlink:href="#g8" y="12716" />
                <use xlink:href="#g10" y="12733" />
                <use xlink:href="#g21" y="12750" />
                <use xlink:href="#g22" y="12767" />
                <use xlink:href="#g23" y="12784" />
                <use xlink:href="#g24" y="12801" />
                <use xlink:href="#g25" y="12818" />
                <use xlink:href="#g26" y="12835" />
                <use xlink:href="#g27" y="12852" />
                <use xlink:href="#g28" y="12869" />
                <use xlink:href="#g29" y="12886" />
                <use xlink:href="#g30" y="12903" />
                <use xlink:href="#g31" y="12920" />
                <use xlink:href="#g32" y="12937" />
                <use xlink:href="#g33" y="12954" />
                <use xlink:href="#g34" y="12971" />
                <use xlink:href="#g41" y="12988" />
                <use xlink:href="#g42" y="13005" />
                <rect x="184" y="13022" width="8" height="17" class="foreground" />
                <use xlink:href="#g45" y="13022" />
            </g>
            <g>
                <use xlink:href="#g8" y="13090" />
                <use xlink:href="#g10" y="13107" />
                <use xlink:href="#g21" y="13124" />
                <use xlink:href="#g22" y="13141" />
                <use xlink:href="#g23" y="13158" />
                <use xlink:href="#g24" y="13175" />
                <use xlink:href="#g25" y="13192" />
                <use xlink:href="#g26" y="13209" />
                <use xlink:href="#g27" y="13226" />
                <use xlink:href="#g28" y="13243" />
                <use xlink:href="#g29" y="13260" />
                <use xlink:href="#g30" y="13277" />
                <use xlink:href="#g31" y="13294" />
                <use xlink:href="#g32" y="13311" />
                <use xlink:href="#g33" y="13328" />
                <use xlink:href="#g34" y="13345" />
                <use xlink:href="#g41" y="13362" />
                <use xlink:href="#g42" y="13379" />
                <rect x="192" y="13396" width="8" height="17" class="foreground" />
                <use xlink:href="#g46" y="13396" />
            </g>
            <g>
                <use xlink:href="#g8" y="13464" />
                <use xlink:href="#g10" y="13481" />
                <use xlink:href="#g21" y="13498" />
                <use xlink:href="#g22" y="13515" />
                <use xlink:href="#g23" y="13532" />
                <use xlink:href="#g24" y="13549" />
                <use xlink:href="#g25" y="13566" />
                <use xlink:href="#g26" y="13583" />
                <use xlink:href="#g27" y="13600" />
                <use xlink:href="#g28" y="13617" />
                <use xlink:href="#g29" y="13634" />
                <use xlink:href="#g30" y="13651" />
                <use xlink:href="#g31" y="13668" />
                <use xlink:href="#g32" y="13685" />
                <use xlink:href="#g33" y="13702" />
                <use xlink:href="#g34" y="13719" />
                <use xlink:href="#g41" y="13736" />
                <use xlink:href="#g42" y="13753" />
                <use xlink:href="#g47" y="13770" />
                <rect x="0" y="13787" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="13787" />
            </g>
            <g>
                <use xlink:href="#g8" y="13838" />
                <use xlink:href="#g10" y="13855" />
                <use xlink:href="#g21" y="13872" />
                <use xlink:href="#g22" y="13889" />
                <use xlink:href="#g23" y="13906" />
                <use xlink:href="#g24" y="13923" />
                <use xlink:href="#g25" y="13940" />
                <use xlink:href="#g26" y="13957" />
                <use xlink:href="#g27" y="13974" />
                <use xlink:href="#g28" y="13991" />
                <use xlink:href="#g29" y="14008" />
                <use xlink:href="#g30" y="14025" />
                <use xlink:href="#g31" y="14042" />
                <use xlink:href="#g32" y="14059" />
                <use xlink:href="#g33" y="14076" />
                <use xlink:href="#g34" y="14093" />
                <use xlink:href="#g41" y="14110" />
                <use xlink:href="#g42" y="14127" />
                <use xlink:href="#g47" y="14144" />
                <use xlink:href="#g48" y="14161" />
                <rect x="0" y="14178" width="8" height="17" class="foreground" />
                <use xlink:href="#g9" y="14178" />
            </g>
        </g>
    </svg>
</svg>
